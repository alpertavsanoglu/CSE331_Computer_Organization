module nor32(a, b, out);
input [31:0] a;
input [31:0] b;
output [31:0] out;

nor nor_0(out[0], b[0], a[0]);
nor nor_1(out[1], b[1], a[1]);
nor nor_2(out[2], b[2], a[2]);
nor nor_3(out[3], b[3], a[3]);
nor nor_4(out[4], b[4], a[4]);
nor nor_5(out[5], b[5], a[5]);
nor nor_6(out[6], b[6], a[6]);
nor nor_7(out[7], b[7], a[7]);
nor nor_8(out[8], b[8], a[8]);
nor nor_9(out[9], b[9], a[9]);
nor nor_10(out[10], b[10], a[10]);
nor nor_11(out[11], b[11], a[11]);
nor nor_12(out[12], b[12], a[12]);
nor nor_13(out[13], b[13], a[13]);
nor nor_14(out[14], b[14], a[14]);
nor nor_15(out[15], b[15], a[15]);
nor nor_16(out[16], b[16], a[16]);
nor nor_17(out[17], b[17], a[17]);
nor nor_18(out[18], b[18], a[18]);
nor nor_19(out[19], b[19], a[19]);
nor nor_20(out[20], b[20], a[20]);
nor nor_21(out[21], b[21], a[21]);
nor nor_22(out[22], b[22], a[22]);
nor nor_23(out[23], b[23], a[23]);
nor nor_24(out[24], b[24], a[24]);
nor nor_25(out[25], b[25], a[25]);
nor nor_26(out[26], b[26], a[26]);
nor nor_27(out[27], b[27], a[27]);
nor nor_28(out[28], b[28], a[28]);
nor nor_29(out[29], b[29], a[29]);
nor nor_30(out[30], b[30], a[30]);
nor nor_31(out[31], b[31], a[31]);


endmodule